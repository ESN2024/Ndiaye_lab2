
module lab2 (
	clk_clk,
	reset_reset_n,
	cnt_3_export,
	cnt_2_export,
	cnt_2_1_export);	

	input		clk_clk;
	input		reset_reset_n;
	input	[7:0]	cnt_3_export;
	input	[7:0]	cnt_2_export;
	input	[7:0]	cnt_2_1_export;
endmodule
